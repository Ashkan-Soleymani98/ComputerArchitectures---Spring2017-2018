module rom(address,data);
input [9:0] address; //needs to be changed
output [31:0] data;	//needs to be changed
reg [31:0] array[1023:0];	//needs to be changed
always @*
begin
// 0.Fetch --> 0
array[0]=32'b0_0001_0010_0_0_00_0010_000_00_0000000000;//0
array[1]=32'b0_0110_0000_0_0_00_1111_001_11_0000000000;//1

// 1.IADD ---> 32
array[32]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//0
array[33]=32'b0_1011_0000_0_0_11_0001_000_00_0000000000;//1
array[34]=32'b0_1101_0000_0_0_00_1111_000_00_0000000000;//2
array[35]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//3
array[36]=32'b0_0000_1100_0_0_00_1111_001_00_0000000000;//4

//	2.ISUB ---> 64
array[64]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//0
array[65]=32'b0_1101_0000_0_0_11_0001_000_00_0000000000;//1
array[66]=32'b0_1011_0000_0_0_00_1111_000_00_0000000000;//2
array[67]=32'b1_0001_1111_0_0_00_1111_000_00_0000000000;//3
array[68]=32'b0_0000_1100_0_0_00_1111_001_00_0000000000;//4

// 3.NOP ---> 96
array[96]=32'b0_1111_1111_0_0_00_1111_001_00_0000000000;//0

// LoadOffset ----> 900
array[900]=32'b0_0001_0010_0_0_00_0010_000_00_0000000000;//0
array[901]=32'b0_1010_0000_0_0_00_0001_000_00_0000000000;//1
array[902]=32'b0_1010_0000_1_0_00_0010_001_10_0000000000;//2

//	Branch ---> 950
array[950]=32'b0_1011_1010_0_0_00_1111_000_00_0000000000;//0
array[951]=32'b0_1101_0010_0_0_00_1111_000_00_0000000000;//1
array[952]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//2
array[953]=32'b0_0010_1100_0_0_00_1111_001_10_0000000000;//3

// 4.GOTO ---> 128
array[128]=32'b0_1111_1111_0_0_00_1111_001_01_1110000100;//0
array[128]=32'b0_1111_1111_0_0_00_1111_001_01_1110110110;//1
array[128]=32'b0_1111_1111_0_0_00_1111_001_00_0000000000;//2

// 5.IFEQ ----> 160
array[160]=32'b0_1111_1111_0_0_00_1111_001_01_1110000100;//0
array[161]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//1
array[162]=32'b0_1011_0000_0_0_00_1111_000_00_0000000000;//2
array[163]=32'b1_0000_1111_0_0_00_1111_000_00_0000000000;//3
array[164]=32'b0_1111_1111_0_0_00_1111_010_01_1110110110;//4
array[165]=32'b0_1111_1111_0_0_00_1111_001_00_0000000000;//5

// 6.IFLT -----> 192
array[192]=32'b0_1111_1111_0_0_00_1111_001_01_1110000100;//0
array[193]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//1
array[194]=32'b0_1011_0000_0_0_00_1111_000_00_0000000000;//2
array[195]=32'b1_0000_1111_0_0_00_1111_000_00_0000000000;//3
array[196]=32'b0_1111_1111_0_0_00_1111_011_01_1110110110;//4
array[197]=32'b0_1111_1111_0_0_00_1111_001_00_0000000000;//5

// 7.IF_ICMPEQ ---> 224 
array[224]=32'b0_1111_1111_0_0_00_1111_001_01_1110000100;//0
array[225]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//1
array[226]=32'b0_1011_0000_0_0_11_0001_000_00_0000000000;//2
array[227]=32'b0_1101_0000_0_0_11_0101_000_00_0000000000;//3
array[228]=32'b0_1111_1111_0_0_00_1111_010_01_1110110110;//4
array[229]=32'b0_1111_1111_0_0_00_1111_001_00_0000000000;//5

//	8.BIPUSH ---> 256
array[256]=32'b0_1111_1111_0_0_00_1111_100_00_0100000101;//0 jmp to 261
array[257]=32'b0_0001_0010_0_0_00_0010_000_00_0000000000;//1
array[258]=32'b0_0111_0000_0_0_01_0101_000_00_0000000000;//2
array[259]=32'b0_0001_0101_0_0_00_1111_000_00_0000000000;//3
array[260]=32'b0_0000_0111_0_0_00_1111_001_00_0000000000;//4
array[261]=32'b0_0001_0101_0_1_00_1111_001_01_1110000100;//5
array[262]=32'b0_0000_1010_0_0_00_1111_001_00_0000000000;//6

// 9.ILOAD ---> 288
array[288]=32'b0_1111_1111_0_0_00_1111_100_00_0100101010;//0 jmp to 298
array[289]=32'b0_0001_0010_0_0_00_0010_000_00_0000000000;//1
array[290]=32'b0_1001_0000_0_0_00_1111_000_00_0000000000;//2
array[291]=32'b0_1011_1001_0_0_00_1111_000_00_0000000000;//3
array[292]=32'b0_1101_0100_0_0_00_1111_000_00_0000000000;//4
array[293]=32'b1_1000_1111_0_0_01_0101_000_00_0000000000;//5
array[294]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//6
array[295]=32'b0_1110_0000_0_0_00_1111_000_00_0000000000;//7
array[296]=32'b0_0001_0101_0_0_00_1111_000_00_0000000000;//8
array[297]=32'b0_0000_1110_0_0_00_1111_001_00_0000000000;//9
array[298]=32'b0_1111_1111_0_1_00_1111_001_01_1110000100;//10
array[299]=32'b0_1011_1010_1_0_00_1111_000_00_0000000000;//11
array[300]=32'b0_1101_0100_0_0_00_1111_000_00_0000000000;//12
array[301]=32'b1_1000_1111_0_0_01_0101_000_00_0000000000;//13
array[302]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//14
array[303]=32'b0_1110_0000_0_0_00_1111_000_00_0000000000;//15
array[304]=32'b0_0001_0101_0_0_00_1111_000_00_0000000000;//16
array[305]=32'b0_0000_1110_0_0_00_1111_001_00_0000000000;//17

//	10.ISTORE ---> 320
array[320]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//0
array[321]=32'b0_1110_0000_0_0_00_1111_100_00_0101001001;//1 jmp to 329
array[322]=32'b0_0001_0010_0_0_00_0010_000_00_0000000000;//2
array[323]=32'b0_1001_0000_0_0_00_1111_000_00_0000000000;//3
array[324]=32'b0_1011_1001_0_0_00_1111_000_00_0000000000;//4
array[325]=32'b0_1101_0100_0_0_00_1111_000_00_0000000000;//5
array[326]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//6
array[327]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//7
array[328]=32'b0_0000_1110_0_0_00_1111_001_00_0000000000;//8
array[329]=32'b0_1111_1111_0_1_00_1111_001_01_1110000100;//9
array[330]=32'b0_1011_1010_1_0_00_1111_000_00_0000000000;//10
array[331]=32'b0_1101_0100_0_0_00_1111_000_00_0000000000;//11
array[332]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//12
array[333]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//13
array[334]=32'b0_0000_1110_0_0_00_1111_001_00_0000000000;//14

//	11.IINC ---> 352
array[352]=32'b0_1111_1111_0_0_00_1111_100_00_0101101100;//0 jmp to 364
array[353]=32'b0_0001_0010_0_0_00_0010_000_00_0000000000;//1
array[354]=32'b0_1001_0000_0_0_00_0001_000_00_0000000000;//2
array[355]=32'b0_1000_0000_0_0_00_0010_000_00_0000000000;//3
array[356]=32'b0_1011_1001_0_0_00_1111_000_00_0000000000;//4
array[357]=32'b0_1101_0100_0_0_00_1111_000_00_0000000000;//5
array[358]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//6
array[359]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//7
array[360]=32'b0_1011_0000_0_0_00_1111_000_00_0000000000;//8
array[361]=32'b0_1101_1000_0_0_00_1111_000_00_0000000000;//9
array[362]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//10
array[363]=32'b0_0000_1100_0_0_00_1111_001_00_0000000000;//11
array[364]=32'b0_1111_1111_0_1_00_1111_001_01_1110000100;//12
array[365]=32'b0_0001_0010_0_0_00_1111_000_00_0000000000;//13
array[366]=32'b0_1000_0000_0_0_00_1111_000_00_0000000000;//14
array[367]=32'b0_1011_1010_1_0_00_1111_000_00_0000000000;//15
array[368]=32'b0_1101_0100_0_0_00_1111_000_00_0000000000;//16
array[369]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//17
array[370]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//18
array[371]=32'b0_1011_0000_0_0_00_1111_000_00_0000000000;//19
array[372]=32'b0_1101_1000_0_0_00_1111_000_00_0000000000;//20
array[373]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//21
array[374]=32'b0_0000_1100_0_0_00_1111_001_00_0000000000;//22

//	12.DUP ---> 384
array[384]=32'b0_0001_0101_0_0_01_0101_000_00_0000000000;//0
array[385]=32'b0_1110_0000_0_0_01_0001_000_00_0000000000;//1
array[386]=32'b0_0000_1110_0_0_00_1111_001_00_0000000000;//2

//	13.IAND ---> 416
array[416]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//0
array[417]=32'b0_1011_0000_0_0_11_0001_000_00_0000000000;//1
array[418]=32'b0_1101_0000_0_0_00_1111_000_00_0000000000;//2
array[419]=32'b1_0111_1111_0_0_00_1111_000_00_0000000000;//3
array[420]=32'b0_0000_1100_0_0_00_1111_001_00_0000000000;//4

// 14.INVOKEVIRTUAL ----> 448
array[448]=32'b0_1111_1111_0_0_00_1111_001_01_1110000100;//0
array[449]=32'b0_1011_1010_1_0_00_1111_000_00_0000000000;//1
array[450]=32'b0_1101_0011_0_0_00_1111_000_00_0000000000;//2
array[451]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//3
array[452]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//4
array[453]=32'b0_0001_0000_0_0_00_1111_000_00_0000000000;//5
array[454]=32'b0_1010_0000_0_0_00_0001_000_00_0000000000;//6
array[455]=32'b0_1010_0000_1_0_00_0001_000_00_0000000000;//7
array[456]=32'b0_1110_0100_0_0_00_1111_000_00_0000000000;//8
array[457]=32'b0_1101_0101_0_0_00_1111_000_00_0000000000;//9
array[458]=32'b0_1011_1010_1_0_00_1111_000_00_0000000000;//10
array[459]=32'b1_0001_1111_0_0_00_1111_000_00_0000000000;//11
array[460]=32'b0_0100_1100_0_0_00_1111_000_00_0000000000;//12
array[461]=32'b0_1010_0000_0_0_00_0001_000_00_0000000000;//13
array[462]=32'b0_1010_0000_1_0_00_0001_000_00_0000000000;//14
array[463]=32'b0_1011_1010_1_0_01_0101_000_00_0000000000;//15
array[464]=32'b0_1101_0101_0_0_01_0100_000_00_0000000000;//16
array[465]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//17
array[466]=32'b0_0101_1100_0_0_00_1111_000_00_0000000000;//18
array[467]=32'b0_0001_0101_0_0_01_0101_000_00_0000000000;//19
array[468]=32'b0_0000_0010_0_0_01_0001_000_00_0000000000;//20
array[469]=32'b0_0000_1110_0_0_00_1111_000_00_0000000000;//21
array[470]=32'b0_0010_0001_0_0_00_1111_001_00_0000000000;//22

//	15.IOR ---> 480
array[480]=32'b0_0001_0101_0_0_11_0101_000_00_0000000000;//0
array[481]=32'b0_1011_0000_0_0_11_0001_000_00_0000000000;//1
array[482]=32'b0_1101_0000_0_0_00_1111_000_00_0000000000;//2
array[483]=32'b1_1001_1111_0_0_00_1111_000_00_0000000000;//3
array[484]=32'b0_0000_1100_0_0_00_1111_001_00_0000000000;//4

// 16.IRETURN ---> 512
array[512]=32'b0_0001_0101_0_0_00_1111_000_00_0000000000;//0
array[513]=32'b0_1110_0000_0_0_11_0001_000_00_0000000000;//1
array[514]=32'b0_0101_0100_0_0_00_1111_000_00_0000000000;//2
array[515]=32'b0_0100_0000_0_0_11_0001_000_00_0000000000;//3
array[516]=32'b0_0010_0000_0_0_00_1111_000_00_0000000000;//4
array[517]=32'b0_0001_0101_0_0_00_1111_000_00_0000000000;//5
array[518]=32'b0_0000_1110_0_0_00_1111_001_00_0000000000;//6

// 17.LDC_W ---> 544
array[544]=32'b0_1111_1111_0_0_00_1111_001_01_1110000100;//0
array[545]=32'b0_1011_1010_1_0_00_1111_000_00_0000000000;//1
array[546]=32'b0_1101_0011_0_0_00_1111_000_00_0000000000;//2
array[547]=32'b1_1000_1111_0_0_00_1111_000_00_0000000000;//3
array[548]=32'b0_0001_1100_0_0_00_1111_000_00_0000000000;//4
array[549]=32'b0_1110_0000_0_0_01_0101_000_00_0000000000;//5
array[550]=32'b0_0001_0101_0_0_00_1111_000_00_0000000000;//6
array[551]=32'b0_0000_1110_0_0_00_1111_001_00_0000000000;//7

//	18.POP ---> 576
array[576]=32'b0_1111_1111_0_0_11_0101_001_00_0000000000;//0

//	19.SWAP ---> 608
array[608]=32'b0_0001_0101_0_0_00_1111_000_00_0000000000;//0
array[609]=32'b0_1110_0000_0_0_11_0001_000_00_0000000000;//1
array[610]=32'b0_1011_0000_0_0_00_1111_000_00_0000000000;//2
array[611]=32'b0_0000_1110_0_0_01_0001_000_00_0000000000;//3
array[612]=32'b0_0000_1011_0_0_00_1111_001_00_0000000000;//4

//	20.WIDE ---> 640
array[640]=32'b0_1111_1111_0_1_00_1111_001_00_0000000000;//0



end
assign data=array[address];
endmodule